module Test (
    output logic led
);
    assign led = 1;

endmodule
