module Layer ();

endmodule
