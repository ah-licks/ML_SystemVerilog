package AF;
    typedef enum {
        Identity,
        Binary_Step,
        ReLU
    } Act_Func;
endpackage
