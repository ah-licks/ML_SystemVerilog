import AF::*;

module Main (
    output logic led
);
    assign led = 1;

endmodule
